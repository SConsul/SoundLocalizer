LPF2 7.95K

.include tl071.txt


*************************************
*Unity Gain HPF cutoff f=10.6Hz

.subckt HPF1 hpf1_IN hpf1_OUT hpf1_COM
x_hpf1   hpf1_1 hpf1_OUT hpf1_3 hpf1_4 hpf1_OUT tl071
vdd_hpf1 hpf1_3 hpf1_COM dc 15 ac 0
vee_hpf1 hpf1_4 hpf1_COM dc -15 ac 0
r_hpf1   hpf1_1 hpf1COM 15k
c_hpf1   hpf1_IN hpf1_1 1u
.ends

*************************************
*Unity Gain LPF cutoff f=7.95kHz
.subckt LPF1 lpf1_IN lpf1_OUT lpf1_COM
x_lpf1   lpf1_COM lpf1_2 lpf1_3 lpf1_4 lpf1_OUT tl071
vdd_lpf1 lpf1_3 lpf1_COM dc 15 ac 0
vee_lpf1 lpf1_4 lpf1_COM dc -15 ac 0
r1_lpf1  lpf1_IN lpf1_2 10k
r2_lpf1  lpf1_2 lpf1_OUT 10k
c_lpf1   lpf1_2 lpf1_OUT 2n
.ends

xh i o 0 HPF1
*xl i o 0 LPF1
vin i 0 dc 0 ac 1

.ac dec 3 100 1Meg
.control
run
plot vdb(o) xlog
.endc
.end
