ZCD
*************************************
*LM111

* CONNECTIONS:
*                POSITIVE INPUT
*                | NEGATIVE INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |  GROUND OR EMITTER OUTPUT
*                | | | | |  |
.SUBCKT LM111_0     3 2 8 4 1 104
*
* PINOUT ORDER +IN -IN V+ V- OUT GND
*----- INPUT STAGE -----
VOS  2 13 DC 0.0007
IEE  8 10 DC 1E-4
RC_Q1  11 4 1517.2
RC_Q2  12 4 1517.2
RE_Q1  10 6 1000
RE_Q2  10 7 1000
Q1  11 3 6 MQ1
Q2  12 13 7 MQ2
*----- SUPPLY CURRENT -----
GSUP  8 4 33 4 1
RSUP  8 45 33333.3
DSUP  45 4 MDS
IIS  4 33 DC 0.00395
RIS  33 4 1 TC=-0.00379747, -3.55271E-20
*----- DELAY VS. OVERDRIVE -----
G1  4 25 12 11 10
RCL  25 4 10
DCL1  25 26 MD0
DCL2  27 25 MD0
VCL1  26 4 DC 9.4
VCL2  4 27 DC 9.4
G2  4 16 25 4 0.01
D3  16 18 MD1
D4  17 16 MD1
V1  18 4 DC 0
V2  4 17 DC 0
*----- INTER STAGE -----
GB  4 20 12 11 100
RB  20 4 10
H1  22 4 POLY(1) V1 0 1089.83 -4491.35
H2  4 21 POLY(1) V2 0 1089.83 -4491.35
DB1  20 22 MDB1
DB2  21 20 MDB1
GT  4 30 20 4 1E-5
RT  30 4 100K
CT  30 4 0.8116E-12
GC  4 35 30 4 0.003448
RC  35 4 1K
*----- OUTPUT SATGE -----
GO  104 40 35 4 -0.01
RO  104 40 10
EOB  41 40 45 4 1
RR  1 104 1MEG
CO  40 104 10P
VOE  42 104 DC -0.0477
QO  1 41 42 MQO
.MODEL MQ1 PNP BF=805.452 XTB=1.1526
.MODEL MQ2 PNP BF=861.069 XTB=1.1526
.MODEL MD0 D IS=1E-10 RS=0.01
.MODEL MD1 D IS=1E-12
.MODEL MDB1 D
.MODEL MDS D IS=1E-16
.MODEL MQO NPN BF=100 RC=13.4286 ISC=1.8E-10
+ BR=10 NR=0.95 CJS=5P CJC=1P TF=2N
.ENDS
.OPTIONS ABSTOL=1P ITL1=150 ITL2=20 ITL4=10 TRTOL=7 

*************************************
*ZCD

Vneg_psd1        14 0 -2.5
Vpos_psd1        13 0 2.5
V1               12 0 sin( 0 1 5K 0 0) 
R2_psd1          13 11 10K 
XU2_psd1         12 0 13 14 11 14 LM111_0

Vneg_psd2        24 0 -2.5
Vpos_psd2        23 0 2.5
V2               22 0 sin( 0 1 5K 0.025m 0) 
R2_psd2          23 21 10K 
XU2_psd2         22 0 23 24 21 24 LM111_0

*************************************
*Half Wave Rectifier_A

.include tl071.txt
.include Diode_1N914.txt

.subckt HWR hwr_IN hwr_OUT hwr_COM
x1 hwr_COM hwr_2 hwr_3 hwr_4 hwr_5 tl071
vdd hwr_3 hwr_COM dc 12 ac 0
vee hwr_4 hwr_COM dc -12 ac 0
r1_hwr hwr_IN hwr_2 10k
d1_hwr hwr_2 hwr_5 1N914
r2_hwr hwr_2 hwr_OUT 10k
d2_hwr hwr_5 hwr_OUT 1N914
*rl 6 0 1k
.ends
*************************************

*xhwr i out 0 HWR

.TEMP 27
.control
tran 2u .6m .2m
plot v(21) - v(11)
.endc
.end
