Family of Curves

.include bfw10.txt

*Usually, the order of terminals are
*drain, gate, source and body respectively

j1 d g gnd bfw10
vgs g gnd dc -2.0 .1V
vds dummy gnd dc 1V
vdummy dummy d dc 0V
.control
*dc vds -.2 0.2 0.01 
dc vgs -2.7 -1.6 0.001 
plot i(vdummy)
.endc
.end

** at vgs swing from -2.8 to 0 Rds varies from 15k to 195

