Narrow Bandpass Filter

.include tl071.txt

x1 1 2 3 4 5 tl071
vdd 3 gnd dc 15 ac 0
vee 4 gnd dc -15 ac 0

r31 2 5 10k
r32 1 gnd 10k
c1 2 6 
r2 6 gnd 
c2 6 5
r1 6 i
vin i gnd ac 1
.ac dec 4 10 1Meg

.control
plot (vdb(5)) xlog
*plot {57.29*vp(5)} xlog
.endc
.end
