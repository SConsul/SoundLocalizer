Integrator

.model ZENER D(bv=2.25v)
.include tl071.txt

.subckt INTEGRATOR IN OUT COM
*   d g s b 
*m1 IN COM s s NMOS4007
*x1 s OUT 3 4 OUT tl071
*vdd 3 COM dc 15 ac 0
*vee 4 COM dc -15 ac 0
r1 IN OUT 1k
c1 OUT COM 1u
vd OUT a dc -0.05
dz a COM ZENER
.ends

vin 1 0 PULSE(-15 15 2ns 2ns 2ns .2ms .2ms)
xint 1 2 0 INTEGRATOR

.control
run
tran 0.01m 4ms 0m
plot v(1) v(2)
.endc
.end
