Inverting Schmitt

.include tl071.txt

x1 1 in 3 4 5 tl071
vdd 3 0 dc 12 ac 0
vee 4 0 dc -12 ac 0
r1 1 0 1k
r2 1 5 1k
vin in 0 dc 1
*vin in 0 sin(0 12 5k 0 0)
.control
*run
*tran 0.001m 1.2ms 0m
dc vin -12 12 0.01
plot v(5) 
.endc
.end
